package core_env_pkg;

  import uvm_pkg::*;
  import bus_resp_agent_pkg::*;

  `include "uvm_macros.svh"
  `include "dv_macros.svh"

  `include "core_env.sv"

endpackage
