package core_test_pkg;

  import uvm_pkg::*;
  import bus_resp_agent_pkg::*;
  import core_env_pkg::*;
  import core_pkg::*;

  `include "uvm_macros.svh"
  `include "dv_macros.svh"

  `include "mem_model.sv"

  `include "core_base_test.sv"
  `include "core_test_lib.sv"

endpackage
