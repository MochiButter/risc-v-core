class core_test_asm extends core_base_test;

endclass
